    Mac OS X            	   2   �                                           ATTR         �   X                  �     com.apple.lastuseddate#PS       �   H  com.apple.macl   ��	`    3�     �Z�ZET�aQ��\��                                                      